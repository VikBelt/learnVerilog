module intro (A,B);

    //define input and output
    input A;
    output B;

    assign B = A;
    
endmodule
